
interface test_if;
   logic [7:0] a;
   logic [7:0] b;
   logic [15:0] prod;


endinterface
