
package vedic_pkg;
   import uvm_pkg::*;

   `include "uvm_macros.svh"
   `include "vedic_env.sv"
endpackage
